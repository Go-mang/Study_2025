module hello_world;
    $display("Hello, World!");
    $finish;

    // git process explanation
    // git init -> initialize git repository
    // git add <file> -> add file to staging area
    // git commit -m "message" -> commit changes, 내가 한 작업에 대한 내용
    // git status -> check status of repository
    // git remote add origin <url> -> add remote repository
    // git push origin master -> push changes to remote repository
    // git pull origin master -> pull changes from remote repository
    
endmodule
