module hello_world;
    $display("Hello, World!");
    $finish;
endmodule
